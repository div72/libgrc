module network

struct AddressBook {
}

pub fn (mut ab AddressBook) modify_trust(ip string, diff int) {}
